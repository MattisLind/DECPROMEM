-- Standard Bipolar 256 x 4 bit PROM 
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity DiagROM is
port(
  address  : in integer range 0 to 1023;
  bitAddress : in integer range 0 to 7;
  data     : out std_logic);
end DiagROM;

architecture logic of DiagROM is
type rom_type is array (0 to 1023) of std_logic_vector(7 downto 0); 
signal dataFromRom: std_logic_vector(7 downto 0);
signal rom : rom_type := ( 

x"1C",x"00",x"FF",x"AA",x"00",x"01",x"04",x"00",x"00",x"00",x"26",x"44",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"1A",x"00",x"00",x"C0",x"02",x"00",x"26",x"10",x"66",x"10",x"A6",x"10",
x"E6",x"10",x"26",x"11",x"66",x"11",x"E6",x"17",x"04",x"00",x"E6",x"17",x"06",x"00",x"E6",x"17",
x"4C",x"00",x"E6",x"17",x"4E",x"00",x"E6",x"11",x"CE",x"65",x"16",x"02",x"9F",x"15",x"04",x"00",
x"DF",x"15",x"E0",x"00",x"06",x"00",x"E6",x"11",x"CE",x"65",x"0E",x"02",x"9F",x"15",x"4C",x"00",
x"DF",x"15",x"E0",x"00",x"4E",x"00",x"37",x"0A",x"7C",x"02",x"F7",x"97",x"C7",x"9F",x"76",x"02",
x"37",x"10",x"6E",x"02",x"17",x"74",x"07",x"00",x"C0",x"65",x"04",x"F8",x"37",x"10",x"5C",x"02",
x"C0",x"65",x"02",x"00",x"37",x"10",x"56",x"02",x"FF",x"35",x"C6",x"00",x"50",x"02",x"03",x"03",
x"F7",x"09",x"F4",x"01",x"01",x"00",x"FF",x"1D",x"4C",x"02",x"40",x"02",x"F7",x"1D",x"46",x"02",
x"42",x"02",x"F7",x"0C",x"3E",x"02",x"F7",x"0C",x"3A",x"02",x"37",x"0A",x"32",x"02",x"FF",x"35",
x"10",x"00",x"2A",x"02",x"03",x"03",x"F7",x"15",x"04",x"00",x"24",x"02",x"F7",x"65",x"04",x"00",
x"1E",x"02",x"FF",x"35",x"20",x"00",x"16",x"02",x"02",x"03",x"F7",x"0C",x"12",x"02",x"C5",x"1D",
x"0E",x"02",x"C5",x"6D",x"10",x"02",x"57",x"21",x"60",x"00",x"29",x"07",x"F7",x"15",x"60",x"00",
x"FE",x"01",x"F7",x"ED",x"00",x"02",x"F8",x"01",x"F7",x"0B",x"F4",x"01",x"03",x"06",x"F7",x"09",
x"96",x"01",x"02",x"00",x"E6",x"11",x"CE",x"65",x"78",x"01",x"9F",x"15",x"04",x"00",x"FF",x"15",
x"01",x"00",x"DA",x"01",x"C0",x"15",x"00",x"20",x"05",x"0A",x"E6",x"15",x"01",x"00",x"E6",x"15",
x"80",x"01",x"05",x"88",x"96",x"25",x"48",x"0A",x"06",x"88",x"C5",x"0B",x"03",x"02",x"F7",x"09",
x"66",x"01",x"03",x"00",x"E6",x"11",x"CE",x"65",x"38",x"01",x"9F",x"15",x"04",x"00",x"E6",x"11",
x"CE",x"65",x"44",x"01",x"9F",x"15",x"4C",x"00",x"FF",x"15",x"07",x"00",x"A0",x"01",x"C3",x"1D",
x"A2",x"01",x"C0",x"15",x"00",x"20",x"C5",x"1F",x"94",x"01",x"C4",x"15",x"01",x"00",x"FF",x"35",
x"20",x"00",x"8A",x"01",x"01",x"03",x"C4",x"0C",x"E6",x"15",x"01",x"00",x"E6",x"10",x"05",x"88",
x"96",x"25",x"C5",x"45",x"40",x"00",x"FF",x"35",x"20",x"00",x"72",x"01",x"0F",x"03",x"FF",x"35",
x"10",x"00",x"68",x"01",x"06",x"02",x"C3",x"35",x"10",x"00",x"08",x"03",x"C5",x"55",x"40",x"00",
x"05",x"01",x"C3",x"35",x"40",x"00",x"02",x"03",x"C5",x"55",x"40",x"00",x"E6",x"1D",x"50",x"01",
x"CE",x"0C",x"83",x"65",x"C5",x"55",x"80",x"00",x"08",x"0A",x"C8",x"0B",x"C5",x"35",x"80",x"00",
x"03",x"03",x"F7",x"09",x"E2",x"00",x"04",x"00",x"C5",x"55",x"80",x"00",x"C8",x"15",x"01",x"01",
x"C8",x"0B",x"C5",x"35",x"80",x"00",x"03",x"03",x"F7",x"09",x"CC",x"00",x"04",x"00",x"06",x"88",
x"35",x"7F",x"FF",x"45",x"04",x"00",x"16",x"01",x"E6",x"11",x"CE",x"65",x"9C",x"00",x"9F",x"15",
x"4C",x"00",x"C1",x"15",x"55",x"55",x"C5",x"15",x"AA",x"AA",x"C3",x"1D",x"06",x"01",x"C4",x"1D",
x"FE",x"00",x"C0",x"15",x"00",x"20",x"E6",x"15",x"04",x"00",x"E6",x"10",x"05",x"88",x"96",x"25",
x"C3",x"65",x"04",x"00",x"C2",x"15",x"00",x"40",x"50",x"10",x"82",x"7E",x"06",x"88",x"0F",x"7F",
x"C4",x"1D",x"DC",x"00",x"C0",x"15",x"00",x"A0",x"C3",x"E5",x"04",x"00",x"E6",x"15",x"04",x"00",
x"E6",x"10",x"05",x"88",x"96",x"25",x"C2",x"15",x"00",x"40",x"60",x"20",x"03",x"02",x"48",x"11",
x"48",x"21",x"03",x"03",x"F7",x"09",x"60",x"00",x"05",x"00",x"89",x"7E",x"06",x"88",x"16",x"7F",
x"C1",x"15",x"01",x"01",x"C4",x"1D",x"A8",x"00",x"C0",x"15",x"00",x"20",x"E6",x"15",x"04",x"00",
x"E6",x"10",x"05",x"88",x"96",x"25",x"C3",x"65",x"04",x"00",x"C2",x"15",x"00",x"40",x"48",x"10",
x"D0",x"0B",x"83",x"7E",x"06",x"88",x"10",x"7F",x"F7",x"09",x"2C",x"00",x"00",x"00",x"96",x"25",
x"F7",x"09",x"24",x"00",x"06",x"00",x"96",x"25",x"F7",x"09",x"1C",x"00",x"07",x"00",x"C5",x"15",
x"01",x"00",x"02",x"00",x"7F",x"21",x"66",x"00",x"04",x"03",x"96",x"25",x"F7",x"09",x"08",x"00",
x"08",x"00",x"C5",x"45",x"80",x"00",x"02",x"00",x"06",x"88",x"3F",x"0A",x"50",x"00",x"FE",x"0B",
x"00",x"00",x"0E",x"02",x"F7",x"6D",x"48",x"00",x"4C",x"00",x"DF",x"9D",x"48",x"00",x"C7",x"9F",
x"E6",x"1D",x"3C",x"00",x"CE",x"00",x"BE",x"65",x"00",x"00",x"FF",x"15",x"01",x"00",x"2E",x"00",
x"C5",x"1D",x"2E",x"00",x"C5",x"0C",x"C5",x"0C",x"05",x"0B",x"B5",x"17",x"EE",x"9F",x"9F",x"15",
x"4E",x"00",x"9F",x"15",x"4C",x"00",x"9F",x"15",x"06",x"00",x"9F",x"15",x"04",x"00",x"85",x"15",
x"84",x"15",x"83",x"15",x"82",x"15",x"81",x"15",x"80",x"15",x"00",x"88",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"39",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DD",x"30"
);

begin

  dataFromRom <= rom(address);
  data <= dataFromRom(7-bitAddress); 
end logic;
